module dec7seg_4bits_hexadec(
    output [6:0] y,    // Saída
    input [3:0] a    // Entrada A
);  

    assign y =  (a == 4'h0) ? 7'b1111110 :
                (a == 4'h1) ? 7'b0110000 :
                (a == 4'h2) ? 7'b1101101 :
                (a == 4'h3) ? 7'b1111001 :
                (a == 4'h4) ? 7'b0110011 :
                (a == 4'h5) ? 7'b1011011 :
                (a == 4'h6) ? 7'b1011111 :
                (a == 4'h7) ? 7'b1110000 :
                (a == 4'h8) ? 7'b1111111 :
                (a == 4'h9) ? 7'b1111011 :
                (a == 4'hA) ? 7'b1110111 :
                (a == 4'hB) ? 7'b0011111 :
                (a == 4'hC) ? 7'b1001110 :
                (a == 4'hD) ? 7'b0111101 :
                (a == 4'hE) ? 7'b1001111 :
                (a == 4'hF) ? 7'b1000111 :
                7'b0000000;
endmodule