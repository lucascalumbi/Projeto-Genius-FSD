
module genius()

endmodule